module memory();

endmodule // memory
module reg_array #(parameter N=16, parameter MSB=16)
	(
      	input clk,
		input we,
		input [$clog2(N)-1:0] addr,
		input [MSB-1:0] data,
      	output [N*MSB-1:0]  data_out 
	);

reg [MSB-1:0] regs [N-1:0];

genvar i;

always @(negedge clk)
begin
if(we)
begin
	regs[addr] <= data;
end
end

generate
	for(i=0;i<N;i=i+1)
	begin
	assign data_out[(i+1)*N-1:N*i] = regs[i];
	end
endgenerate





endmodule // input_regs
module top
(
input CLK,
		);